-- Testbench de Decimal a display 7 segmentos de las decenas
library IEEE;
use IEEE.std_logic_1164.all;

entity tb_of_bcd7seg_dec is
end entity;

architecture tb of tb_of_bcd7seg_dec is
component bcd7seg_dec is
Port ( 
        decenas: integer range 0 to 9;
        segmentos_dec : out std_logic_vector (6 downto 0)
);
end component;

signal decenas_IN : integer;
signal segmentos_dec_OUT : std_logic_vector (6 downto 0);

begin

UUT : bcd7seg_dec port map (
	decenas => decenas_IN,
    segmentos_dec => segmentos_dec_OUT
);


stimulation_signals : process
begin

decenas_IN <= 9;
wait for 5 ns;
decenas_IN <= 8;
wait for 20ns;
decenas_IN <= 7;
wait for 5 ns;
decenas_IN <= 6;
wait for 15 ns;
decenas_IN <= 5;
wait for 5 ns;
decenas_IN <= 4;
wait for 10 ns;
decenas_IN <= 3;
wait for 5 ns;
decenas_IN <= 2;
wait for 15 ns;
decenas_IN <= 1;
wait for 5 ns;
decenas_IN <= 0;
wait for 10 ns;
-- Run Time:100 ns
	
end process;


end tb;